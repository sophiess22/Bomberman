5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 
5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 
5'hB, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 
5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA
potion:
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h3, 5'h3, 5'h3, 5'h3, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h3, 5'h3, 5'h3, 5'h3, 5'hE, 5'hE, 5'hE, 5'hE, 5'h3, 5'h3, 5'h3, 5'h3, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hC, 5'hB, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hC, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'hC, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hA, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hC, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hA, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hC, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hA, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h
shoe:
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h3, 5'h3, 5'h3, 5'h3, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'h1, 5'hC, 5'hC, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h0, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h1, 5'h1, 5'h1, 5'h1, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'hC, 5'hC, 5'hC, 5'h0, 5'hA, 5'hB, 5'hB, 5'hA, 5'hA, 5'hC, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'h0, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hA, 5'hA, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'h0, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'h0, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hC, 5'hC, 5'hC, 5'hC, 5'h0, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'hA, 5'hB, 5'hB, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hC, 5'hB, 5'hC, 5'h0, 5'hC, 5'hC, 5'hB, 5'hB, 5'hB, 5'hC, 5'hC, 5'hA, 5'hA, 5'h0, 5'hA, 5'hA, 5'hA, 5'h0, 5'h0, 5'h8, 5'hB, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'hC, 5'hB, 5'hB, 5'hC, 5'hC, 5'hC, 5'hB, 5'hB, 5'hC, 5'hC, 5'hB, 5'hA, 5'hA, 5'hA, 5'hA, 5'hB, 5'hA, 5'hA, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hA, 5'hA, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'hB, 5'hB, 5'hB, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h0, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'h8, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 
5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF, 5'hF


0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 
0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0